grammar edu:umn:cs:melt:exts:ableC:interval;

exports edu:umn:cs:melt:exts:ableC:interval:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:interval:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:string;