grammar edu:umn:cs:melt:exts:ableC:interval:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:interval:concretesyntax:typeExpr;
exports edu:umn:cs:melt:exts:ableC:interval:concretesyntax:constructor;